`timescale 1ns / 1ps

module tb_imit_signal(

    );
endmodule
